library verilog;
use verilog.vl_types.all;
entity CPUProject_vlg_vec_tst is
end CPUProject_vlg_vec_tst;
