module ALU_TB ();



endmodule